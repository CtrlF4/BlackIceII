// Test verilog file for atom


module testand(a, b, f);
  input a,b;
  output f;

  assign f = a + b;


endmoudle testand:
